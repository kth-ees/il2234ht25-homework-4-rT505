module constraint_random_tb;

//write your code here

endmodule


