module imc_tb;

// Testbench code goes here
endmodule