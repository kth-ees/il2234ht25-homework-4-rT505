module input_out_wrapper_tb;
// Testbench code goes here
endmodule