module iab_tb;

// Testbench code goes here
endmodule